module  decoder3_8(
        input         [ 2: 0]  a                        ,//输入端口a,[2:0]表示位宽
        input                  g1                       ,//使能信号1
        input                  g2                       ,//使能信号2
        input                  g3                       ,//使能信号3
        output  reg   [ 7: 0]  y                         //输出端口y，[7:0]表示位宽
);
//=====================================================================\
// ********** Define Parameter and Internal Signals *************
//=====================================================================/




//======================================================================
// ***************      Main    Code    ****************
//======================================================================
always  @(*) begin
        if({g3,g2,g1} != 3'b001) //g3,g2,g1位使能信号，当他们为001是使能
           y        <=      8'h00;
        else 
           case(a)
              3'b000:   y       <=      8'b0000_0001; 
              3'b001:   y       <=      8'b0000_0010; 
              3'b010:   y       <=      8'b0000_0100; 
              3'b011:   y       <=      8'b0000_1000; 
              3'b100:   y       <=      8'b0001_0000; 
              3'b101:   y       <=      8'b0010_0000; 
              3'b110:   y       <=      8'b0100_0000; 
              3'b111:   y       <=      8'b1000_0000; 
           endcase
end





endmodule
